package my_testbench_pkg;
  import uvm_pkg::*;

  `include "memory_pkt.sv"
  `include "memory_coverage.sv"
  `include "memory_scoreboard.sv"
  `include "memory_monitor.sv"
  `include "memory_sequencer.sv"
  `include "memory_traffic_sequence.sv"
  `include "memory_driver.sv"
  `include "memory_agent.sv"
  `include "memory_env.sv"
  `include "my_test.sv"

endpackage